module ALU();
    // TODO
endmodule