`define OP_SPECIAL  6'b000000
`define FN_ADD      6'b100000
`define FN_ADDU     6'b100001
`define FN_AND      6'b100100
`define FN_BREAK    6'b001101
`define FN_DIV      6'b011010
`define FN_DIVU     6'b011011
`define FN_JR       6'b001000
`define FN_MFHI     6'b010000
`define FN_MFLO     6'b010010
`define FN_MTHI     6'b010001
`define FN_MTLO     6'b010011
`define FN_MULT     6'b011000
`define FN_MULTU    6'b011001
`define FN_NOR      6'b100111
`define FN_OR       6'b100101
`define FN_SLL      6'b000000
`define FN_SLLV     6'b000100
`define FN_SLT      6'b101010
`define FN_SLTU     6'b101011
`define FN_SRA      6'b000011
`define FN_SRAV     6'b000111
`define FN_SRL      6'b000010
`define FN_SRLV     6'b000110
`define FN_SUB      6'b100010
`define FN_SUBU     6'b100011
`define FN_SYSCALL  6'b001100
`define FN_XOR      6'b100110

`define OP_ADDI     6'b001000
`define OP_ADDIU    6'b001001
`define OP_ANDI     6'b001100
`define OP_LB       6'b100000
`define OP_LBU      6'b100100
`define OP_LH       6'b100001
`define OP_LHU      6'b100101
`define OP_LUI      6'b001111
`define OP_LW       6'b100011
`define OP_LWL      6'b100010
`define OP_LWR      6'b100110
`define OP_ORI      6'b001101
`define OP_SB       6'b101000
`define OP_SH       6'b101001
`define OP_SLTI     6'b001010
`define OP_SLTIU    6'b001011
`define OP_SW       6'b101011
`define OP_SWL      6'b101010
`define OP_SWR      6'b101110
`define OP_XORI     6'b001110
`define OP_BEQ      6'b000100
`define OP_REGIMM   6'b000001
`define OP_BGTZ     6'b000111
`define OP_BLEZ     6'b000110
`define OP_BNE      6'b000101
`define OP_J        6'b000010
`define OP_JAL      6'b000011
`define OP_JALR     6'b001001

`define REGIMM_BGEZ     5'b00001
`define REGIMM_BGEZAL   5'b10001
`define REGIMM_BLTZ     5'b00000
`define REGIMM_BLTZAL   5'b10000