module PC();
    // TODO
endmodule